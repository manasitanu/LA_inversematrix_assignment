`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
//Student: Manasi Dubey
// 
// Create Date:    10:13:39 10/07/2016 
// Design Name: 
// Module Name:    matrix_inverse 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module matrix_inverse(clk);

input clk;
real a[0:4][0:9];

always@(posedge clk)
begin
		//initialising the inputs
		a[0][0]=16'd1;
		a[0][1]=16'd2;
		a[0][2]=16'd1;
		a[0][3]=16'd0;
		a[0][4]=16'd0;
		a[0][5]=16'd1;
		a[0][6]=16'd0;
		a[0][7]=16'd0;
		a[0][8]=16'd0;
		a[0][9]=16'd0;
		
		a[1][0]=16'd0;
	   a[1][1]=16'd1;
      a[1][2]=16'd2;
      a[1][3]=16'd1;
      a[1][4]=16'd0;
		a[1][5]=16'd0;
		a[1][6]=16'd1;
		a[1][7]=16'd0;
		a[1][8]=16'd0;
		a[1][9]=16'd0;

		a[2][0]=16'd0;
      a[2][1]=16'd0;
		a[2][2]=16'd1;
		a[2][3]=16'd2;
		a[2][4]=16'd1;
		a[2][5]=16'd0;
		a[2][6]=16'd0;
		a[2][7]=16'd1;
		a[2][8]=16'd0;
		a[2][9]=16'd0;
		
		
		a[3][0]=16'd0;
		a[3][1]=16'd0;
		a[3][2]=16'd0;
		a[3][3]=16'd1;
		a[3][4]=16'd2;
		a[3][5]=16'd0;
		a[3][6]=16'd0;
		a[3][7]=16'd0;
		a[3][8]=16'd1;
		a[3][9]=16'd0;
		
		a[4][0]=16'd0;
		a[4][1]=16'd0;
		a[4][2]=16'd0;
		a[4][3]=16'd0;
		a[4][4]=16'd1;
		a[4][5]=16'd0;
		a[4][6]=16'd0;
		a[4][7]=16'd0;
		a[4][8]=16'd0;
		a[4][9]=16'd1;


		//if first element is not equal to zero then perform the task of addition or subtraction or scalar multiplication
		if(a[0][0]!=0)
		begin
		//making first element equals to 1
		a[0][0]=a[0][0]/a[0][0];
		a[0][1]=a[0][1]/a[0][0];
		a[0][2]=a[0][2]/a[0][0];
		a[0][3]=a[0][3]/a[0][0];
		a[0][4]=a[0][4]/a[0][0];
		a[0][5]=a[0][5]/a[0][0];
		a[0][6]=a[0][6]/a[0][0];
		a[0][7]=a[0][7]/a[0][0];
		a[0][8]=a[0][8]/a[0][0];
		a[0][9]=a[0][9]/a[0][0];
		
		//making element at a[1][0] equals to 0
		a[1][0]=a[1][0]+(-a[1][0]*a[0][0]);
		a[1][1]=a[1][1]+(-a[1][0]*a[0][1]);
		a[1][2]=a[1][2]+(-a[1][0]*a[0][2]);
		a[1][3]=a[1][3]+(-a[1][0]*a[0][3]);
		a[1][4]=a[1][4]+(-a[1][0]*a[0][4]);
		a[1][5]=a[1][5]+(-a[1][0]*a[0][5]);
		a[1][6]=a[1][6]+(-a[1][0]*a[0][6]);
		a[1][7]=a[1][7]+(-a[1][0]*a[0][7]);
		a[1][8]=a[1][8]+(-a[1][0]*a[0][8]);
		a[1][9]=a[1][9]+(-a[1][0]*a[0][9]);
		
		
		
		//making element at a[2][0] equals to 0
		a[2][0]=a[2][0]+(-a[2][0]*a[0][0]);
		a[2][1]=a[2][1]+(-a[2][0]*a[0][1]);
		a[2][2]=a[2][2]+(-a[2][0]*a[0][2]);
		a[2][3]=a[2][3]+(-a[2][0]*a[0][3]);
		a[2][4]=a[2][4]+(-a[2][0]*a[0][4]);
		a[2][5]=a[2][5]+(-a[2][0]*a[0][5]);
		a[2][6]=a[2][6]+(-a[2][0]*a[0][6]);
		a[2][7]=a[2][7]+(-a[2][0]*a[0][7]);
		a[2][8]=a[2][8]+(-a[2][0]*a[0][8]);
		a[2][9]=a[2][9]+(-a[2][0]*a[0][9]);
		
				
		//making element at a[3][0] equals to 0
		a[3][0]=a[3][0]+(-a[3][0]*a[0][0]);
		a[3][1]=a[3][1]+(-a[3][0]*a[0][1]);
		a[3][2]=a[3][2]+(-a[3][0]*a[0][2]);
		a[3][3]=a[3][3]+(-a[3][0]*a[0][3]);
		a[3][4]=a[3][4]+(-a[3][0]*a[0][4]);
		a[3][5]=a[3][5]+(-a[3][0]*a[0][5]);
		a[3][6]=a[3][6]+(-a[3][0]*a[0][6]);
		a[3][7]=a[3][7]+(-a[3][0]*a[0][7]);
		a[3][8]=a[3][8]+(-a[3][0]*a[0][8]);
		a[3][9]=a[3][9]+(-a[3][0]*a[0][9]);

				
		//making element at a[4][0] equals to 0
		a[4][0]=a[4][0]+(-a[4][0]*a[0][0]);
		a[4][1]=a[4][1]+(-a[4][0]*a[0][1]);
		a[4][2]=a[4][2]+(-a[4][0]*a[0][2]);
		a[4][3]=a[4][3]+(-a[4][0]*a[0][3]);
		a[4][4]=a[4][4]+(-a[4][0]*a[0][4]);
		a[4][5]=a[4][5]+(-a[4][0]*a[0][5]);
		a[4][6]=a[4][6]+(-a[4][0]*a[0][6]);
		a[4][7]=a[4][7]+(-a[4][0]*a[0][7]);
		a[4][8]=a[4][8]+(-a[4][0]*a[0][8]);
		a[4][9]=a[4][9]+(-a[4][0]*a[0][9]);

		end
		
		//making element at a[1][1] equals to 1
		if(a[1][1]!=0)
		begin
		a[1][0]=a[1][0]/a[1][1];
		a[1][1]=a[1][1]/a[1][1];
		a[1][2]=a[1][2]/a[1][1];
		a[1][3]=a[1][3]/a[1][1];
		a[1][4]=a[1][4]/a[1][1];
		a[1][5]=a[1][5]/a[1][1];
		a[1][6]=a[1][6]/a[1][1];
		a[1][7]=a[1][7]/a[1][1];
		a[1][8]=a[1][8]/a[1][1];
		a[1][9]=a[1][9]/a[1][1];
		
		//making element at a[2][1] equals to 0
		a[2][0]=a[2][0]+(-a[2][1]*a[1][0]);
		a[2][1]=a[2][1]+(-a[2][1]*a[1][1]);
		a[2][2]=a[2][2]+(-a[2][1]*a[1][2]);
		a[2][3]=a[2][3]+(-a[2][1]*a[1][3]);
		a[2][4]=a[2][4]+(-a[2][1]*a[1][4]);
		a[2][5]=a[2][5]+(-a[2][1]*a[1][5]);
		a[2][6]=a[2][6]+(-a[2][1]*a[1][6]);
		a[2][7]=a[2][7]+(-a[2][1]*a[1][7]);
		a[2][8]=a[2][8]+(-a[2][1]*a[1][8]);
		a[2][9]=a[2][9]+(-a[2][1]*a[1][9]);
		
		//making element at a[3][1] equals to 0
		a[3][0]=a[3][0]+(-a[3][1]*a[1][0]);
		a[3][1]=a[3][1]+(-a[3][1]*a[1][1]);
		a[3][2]=a[3][2]+(-a[3][1]*a[1][2]);
		a[3][3]=a[3][3]+(-a[3][1]*a[1][3]);
		a[3][4]=a[3][4]+(-a[3][1]*a[1][4]);
		a[3][5]=a[3][5]+(-a[3][1]*a[1][5]);
		a[3][6]=a[3][6]+(-a[3][1]*a[1][6]);
		a[3][7]=a[3][7]+(-a[3][1]*a[1][7]);
		a[3][8]=a[3][8]+(-a[3][1]*a[1][8]);
		a[3][9]=a[3][9]+(-a[3][1]*a[1][9]);
	
		//making element at a[4][1] equals to 0
		a[4][0]=a[4][0]+(-a[4][1]*a[1][0]);
		a[4][1]=a[4][1]+(-a[4][1]*a[1][1]);
		a[4][2]=a[4][2]+(-a[4][1]*a[1][2]);
		a[4][3]=a[4][3]+(-a[4][1]*a[1][3]);
		a[4][4]=a[4][4]+(-a[4][1]*a[1][4]);
		a[4][5]=a[4][5]+(-a[4][1]*a[1][5]);
		a[4][6]=a[4][6]+(-a[4][1]*a[1][6]);
		a[4][7]=a[4][7]+(-a[4][1]*a[1][7]);
		a[4][8]=a[4][8]+(-a[4][1]*a[1][8]);
		a[4][9]=a[4][9]+(-a[4][1]*a[1][9]);
		end
		
		//making element at a[2][2] equals to 1
		if(a[2][2]!=0)
		begin
		a[2][0]=a[2][0]/a[2][2];
		a[2][1]=a[2][1]/a[2][2];
		a[2][2]=a[2][2]/a[2][2];
		a[2][3]=a[2][3]/a[2][2];
		a[2][4]=a[2][4]/a[2][2];
		a[2][5]=a[2][5]/a[2][2];
		a[2][6]=a[2][6]/a[2][2];
		a[2][7]=a[2][7]/a[2][2];
		a[2][8]=a[2][8]/a[2][2];
		a[2][9]=a[2][9]/a[2][2];
		
		//making element at a[3][2] equals to 0
		a[3][0]=a[3][0]+(-a[3][2]*a[2][0]);
		a[3][1]=a[3][1]+(-a[3][2]*a[2][1]);
		a[3][2]=a[3][2]+(-a[3][2]*a[2][2]);
		a[3][3]=a[3][3]+(-a[3][2]*a[2][3]);
		a[3][4]=a[3][4]+(-a[3][2]*a[2][4]);
		a[3][5]=a[3][5]+(-a[3][2]*a[2][5]);
		a[3][6]=a[3][6]+(-a[3][2]*a[2][6]);
		a[3][7]=a[3][7]+(-a[3][2]*a[2][7]);
		a[3][8]=a[3][8]+(-a[3][2]*a[2][8]);
		a[3][9]=a[3][9]+(-a[3][2]*a[2][9]);

		//making element at a[3][3] equals to 0
		a[4][0]=a[4][0]+(-a[4][2]*a[2][0]);
		a[4][1]=a[4][1]+(-a[4][2]*a[2][1]);
		a[4][2]=a[4][2]+(-a[4][2]*a[2][2]);
		a[4][3]=a[4][3]+(-a[4][2]*a[2][3]);
		a[4][4]=a[4][4]+(-a[4][2]*a[2][4]);
		a[4][5]=a[4][5]+(-a[4][2]*a[2][5]);
		a[4][6]=a[4][6]+(-a[4][2]*a[2][6]);
		a[4][7]=a[4][7]+(-a[4][2]*a[2][7]);
		a[4][8]=a[4][8]+(-a[4][2]*a[2][8]);
		a[4][9]=a[4][9]+(-a[4][2]*a[2][9]);
		end
		
		//making element at a[3][3] equals to 1
		if(a[3][3]!=0)
		begin
		a[3][0]=a[3][0]/a[3][3];
		a[3][1]=a[3][1]/a[3][3];
		a[3][2]=a[3][2]/a[3][3];
		a[3][3]=a[3][3]/a[3][3];
		a[3][4]=a[3][4]/a[3][3];
		a[3][5]=a[3][5]/a[3][3];
		a[3][6]=a[3][6]/a[3][3];
		a[3][7]=a[3][7]/a[3][3];
		a[3][8]=a[3][8]/a[3][3];
		a[3][9]=a[3][9]/a[3][3];

		//making element at a[4][3] equals to 0
		a[4][0]=a[4][0]+(-a[4][3]*a[3][0]);
		a[4][1]=a[4][1]+(-a[4][3]*a[3][1]);
		a[4][2]=a[4][2]+(-a[4][3]*a[3][2]);
		a[4][3]=a[4][3]+(-a[4][3]*a[3][3]);
		a[4][4]=a[4][4]+(-a[4][3]*a[3][4]);
		a[4][5]=a[4][5]+(-a[4][3]*a[3][5]);
		a[4][6]=a[4][6]+(-a[4][3]*a[3][6]);
		a[4][7]=a[4][7]+(-a[4][3]*a[3][7]);
		a[4][8]=a[4][8]+(-a[4][3]*a[3][8]);
		a[4][9]=a[4][9]+(-a[4][3]*a[3][9]);
		end
		
		//making element at a[4][4] equals to 1
		if(a[4][4]!=0)
		begin
		a[4][0]=a[4][0]/a[4][4];
		a[4][1]=a[4][1]/a[4][4];
		a[4][2]=a[4][2]/a[4][4];
		a[4][3]=a[4][3]/a[4][4];
		a[4][4]=a[4][4]/a[4][4];
		a[4][5]=a[4][5]/a[4][4];
		a[4][6]=a[4][6]/a[4][4];
		a[4][7]=a[4][7]/a[4][4];
		a[4][8]=a[4][8]/a[4][4];
		a[4][9]=a[4][9]/a[4][4];
		end
		
		
		//making element at a[0][1] equals to 0
		a[0][0]=a[0][0]+(-a[0][1]*a[1][0]);
		a[0][1]=a[0][1]+(-a[0][1]*a[1][1]);
		a[0][2]=a[0][2]+(-a[0][1]*a[1][2]);
		a[0][3]=a[0][3]+(-a[0][1]*a[1][3]);
		a[0][4]=a[0][4]+(-a[0][1]*a[1][4]);
		a[0][5]=a[0][5]+(-a[0][1]*a[1][5]);
		a[0][6]=a[0][6]+(-a[0][1]*a[1][6]);
		a[0][7]=a[0][7]+(-a[0][1]*a[1][7]);
		a[0][8]=a[0][8]+(-a[0][1]*a[1][8]);
		a[0][9]=a[0][9]+(-a[0][1]*a[1][9]);
		
		//making element at a[1][2] equals to 0
		a[1][0]=a[1][0]+(-a[1][2]*a[2][0]);
		a[1][1]=a[1][1]+(-a[1][2]*a[2][1]);
		a[1][2]=a[1][2]+(-a[1][2]*a[2][2]);
		a[1][3]=a[1][3]+(-a[1][2]*a[2][3]);
		a[1][4]=a[1][4]+(-a[1][2]*a[2][4]);
		a[1][5]=a[1][5]+(-a[1][2]*a[2][5]);
		a[1][6]=a[1][6]+(-a[1][2]*a[2][6]);
		a[1][7]=a[1][7]+(-a[1][2]*a[2][7]);
		a[1][8]=a[1][8]+(-a[1][2]*a[2][8]);
		a[1][9]=a[1][9]+(-a[1][2]*a[2][9]);
		
		//making element at a[0][2] equals to 0
		a[0][0]=a[0][0]+(-a[0][2]*a[2][0]);
		a[0][1]=a[0][1]+(-a[0][2]*a[2][1]);
		a[0][2]=a[0][2]+(-a[0][2]*a[2][2]);
		a[0][3]=a[0][3]+(-a[0][2]*a[2][3]);
		a[0][4]=a[0][4]+(-a[0][2]*a[2][4]);
		a[0][5]=a[0][5]+(-a[0][2]*a[2][5]);
		a[0][6]=a[0][6]+(-a[0][2]*a[2][6]);
		a[0][7]=a[0][7]+(-a[0][2]*a[2][7]);
		a[0][8]=a[0][8]+(-a[0][2]*a[2][8]);
		a[0][9]=a[0][9]+(-a[0][2]*a[2][9]);
		
		//making element at a[0][3] equals to 0
		a[0][0]=a[0][0]+(-a[0][3]*a[3][0]);
		a[0][1]=a[0][1]+(-a[0][3]*a[3][1]);
		a[0][2]=a[0][2]+(-a[0][3]*a[3][2]);
		a[0][3]=a[0][3]+(-a[0][3]*a[3][3]);
		a[0][4]=a[0][4]+(-a[0][3]*a[3][4]);
		a[0][5]=a[0][5]+(-a[0][3]*a[3][5]);
		a[0][6]=a[0][6]+(-a[0][3]*a[3][6]);
		a[0][7]=a[0][7]+(-a[0][3]*a[3][7]);
		a[0][8]=a[0][8]+(-a[0][3]*a[3][8]);
		a[0][9]=a[0][9]+(-a[0][3]*a[3][9]);
		
		//making element at a[1][3] equals to 0
		a[1][0]=a[1][0]+(-a[1][3]*a[3][0]);
		a[1][1]=a[1][1]+(-a[1][3]*a[3][1]);
		a[1][2]=a[1][2]+(-a[1][3]*a[3][2]);
		a[1][3]=a[1][3]+(-a[1][3]*a[3][3]);
		a[1][4]=a[1][4]+(-a[1][3]*a[3][4]);
		a[1][5]=a[1][5]+(-a[1][3]*a[3][5]);
		a[1][6]=a[1][6]+(-a[1][3]*a[3][6]);
		a[1][7]=a[1][7]+(-a[1][3]*a[3][7]);
		a[1][8]=a[1][8]+(-a[1][3]*a[3][8]);
		a[1][9]=a[1][9]+(-a[1][3]*a[3][9]);
		
		//making element at a[2][3] equals to 0
		a[2][0]=a[2][0]+(-a[2][3]*a[3][0]);
		a[2][1]=a[2][1]+(-a[2][3]*a[3][1]);
		a[2][2]=a[2][2]+(-a[2][3]*a[3][2]);
		a[2][3]=a[2][3]+(-a[2][3]*a[3][3]);
		a[2][4]=a[2][4]+(-a[2][3]*a[3][4]);
		a[2][5]=a[2][5]+(-a[2][3]*a[3][5]);
		a[2][6]=a[2][6]+(-a[2][3]*a[3][6]);
		a[2][7]=a[2][7]+(-a[2][3]*a[3][7]);
		a[2][8]=a[2][8]+(-a[2][3]*a[3][8]);
		a[2][9]=a[2][9]+(-a[2][3]*a[3][9]);
		
		
		//making element at a[0][4] equals to 0
		a[0][0]=a[0][0]+(-a[0][4]*a[4][0]);
		a[0][1]=a[0][1]+(-a[0][4]*a[4][1]);
		a[0][2]=a[0][2]+(-a[0][4]*a[4][2]);
		a[0][3]=a[0][3]+(-a[0][4]*a[4][3]);
		a[0][4]=a[0][4]+(-a[0][4]*a[4][4]);
		a[0][5]=a[0][5]+(-a[0][4]*a[4][5]);
		a[0][6]=a[0][6]+(-a[0][4]*a[4][6]);
		a[0][7]=a[0][7]+(-a[0][4]*a[4][7]);
		a[0][8]=a[0][8]+(-a[0][4]*a[4][8]);
		a[0][9]=a[0][9]+(-a[0][4]*a[4][9]);
		
		//making element at a[1][4] equals to 0
		a[1][0]=a[1][0]+(-a[1][4]*a[4][0]);
		a[1][1]=a[1][1]+(-a[1][4]*a[4][1]);
		a[1][2]=a[1][2]+(-a[1][4]*a[4][2]);
		a[1][3]=a[1][3]+(-a[1][4]*a[4][3]);
		a[1][4]=a[1][4]+(-a[1][4]*a[4][4]);
		a[1][5]=a[1][5]+(-a[1][4]*a[4][5]);
		a[1][6]=a[1][6]+(-a[1][4]*a[4][6]);
		a[1][7]=a[1][7]+(-a[1][4]*a[4][7]);
		a[1][8]=a[1][8]+(-a[1][4]*a[4][8]);
		a[1][9]=a[1][9]+(-a[1][4]*a[4][9]);
		
		//making element at a[2][34] equals to 0
		a[2][0]=a[2][0]+(-a[2][4]*a[4][0]);
		a[2][1]=a[2][1]+(-a[2][4]*a[4][1]);
		a[2][2]=a[2][2]+(-a[2][4]*a[4][2]);
		a[2][3]=a[2][3]+(-a[2][4]*a[4][3]);
		a[2][4]=a[2][4]+(-a[2][4]*a[4][4]);
		a[2][5]=a[2][5]+(-a[2][4]*a[4][5]);
		a[2][6]=a[2][6]+(-a[2][4]*a[4][6]);
		a[2][7]=a[2][7]+(-a[2][4]*a[4][7]);
		a[2][8]=a[2][8]+(-a[2][4]*a[4][8]);
		a[2][9]=a[2][9]+(-a[2][4]*a[4][9]);
		
		//making element at a[3][4] equals to 0
		a[3][0]=a[3][0]+(-a[3][4]*a[4][0]);
		a[3][1]=a[3][1]+(-a[3][4]*a[4][1]);
		a[3][2]=a[3][2]+(-a[3][4]*a[4][2]);
		a[3][3]=a[3][3]+(-a[3][4]*a[4][3]);
		a[3][4]=a[3][4]+(-a[3][4]*a[4][4]);
		a[3][5]=a[3][5]+(-a[3][4]*a[4][5]);
		a[3][6]=a[3][6]+(-a[3][4]*a[4][6]);
		a[3][7]=a[3][7]+(-a[3][4]*a[4][7]);
		a[3][8]=a[3][8]+(-a[3][4]*a[4][8]);
		a[3][9]=a[3][9]+(-a[3][4]*a[4][9]);
		

		//to display the output
		$write("%f	",a[0][5]);
		$write("%f	",a[0][6]);
		$write("%f	",a[0][7]);
		$write("%f	",a[0][8]);
		$display("%f",a[0][9]);
		
		$write("%f	",a[1][5]);
		$write("%f	",a[1][6]);
		$write("%f	",a[1][7]);
		$write("%f	",a[1][8]);
		$display("%f",a[1][9]);
		
		$write("%f	",a[2][5]);
		$write("%f	",a[2][6]);
		$write("%f	",a[2][7]);
		$write("%f	",a[2][8]);
		$display("%f",a[2][9]);
		
		$write("%f	",a[3][5]);
		$write("%f	",a[3][6]);
		$write("%f	",a[3][7]);
		$write("%f	",a[3][8]);
		$display("%f",a[3][9]);
		
		$write("%f	",a[4][5]);
		$write("%f	",a[4][6]);
		$write("%f	",a[4][7]);
		$write("%f	",a[4][8]);
		$display("%f",a[4][9]);

		
		
end

endmodule
